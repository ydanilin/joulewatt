** Profile: "SCHEMATIC1-Voltref"  [ C:\USERS\YURETZZ\DOCUMENTS\������ �����������\�������������\VAHDIODIKA\CHAPTER01\PSPICE\Voltref02\voltref02-pspicefiles\schematic1\voltref.sim ] 

** Creating circuit file "Voltref.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../voltref02-pspicefiles/voltref02.lib" 
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 
.stmlib "C:\Cadence\SPB_16.3\tools\pspice\library\nom.lib" 

*Analysis directives: 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
