** Profile: "SCHEMATIC1-Res_sweep"  [ C:\USERS\YURETZZ\DOCUMENTS\������ �����������\�������������\VAHDIODIKA\CHAPTER01\PSPICE\Voltref02\Voltref02-PSpiceFiles\SCHEMATIC1\Res_sweep.sim ] 

** Creating circuit file "Res_sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../voltref02-pspicefiles/voltref02.lib" 
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 
.stmlib "C:\Cadence\SPB_16.3\tools\pspice\library\nom.lib" 

*Analysis directives: 
.DC LIN PARAM rvariable 60 140 0.001 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
