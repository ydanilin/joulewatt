** Profile: "SCHEMATIC1-Vah-bias"  [ C:\USERS\YURETZZ\DOCUMENTS\������ �����������\�������������\VAHDIODIKA\CHAPTER01\PSPICE\Vah02\Two-diodikas-PSpiceFiles\SCHEMATIC1\Vah-bias.sim ] 

** Creating circuit file "Vah-bias.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../two-diodikas-pspicefiles/two-diodikas.lib" 
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 
.stmlib "C:\Cadence\SPB_16.3\tools\pspice\library\nom.lib" 

*Analysis directives: 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
