** Profile: "SCHEMATIC1-Vreference"  [ C:\USERS\YURETZZ\DOCUMENTS\������ �����������\�������������\VAHDIODIKA\CHAPTER01\PSPICE\Voltref01\Voltref-PSpiceFiles\SCHEMATIC1\Vreference.sim ] 

** Creating circuit file "Vreference.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 
.stmlib "C:\Cadence\SPB_16.3\tools\pspice\library\nom.lib" 

*Analysis directives: 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
